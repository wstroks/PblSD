`ifndef ALUOP
`define ALUOP

`define ALU_ADDU 5'd0
`define ALU_ADD  5'd1
`define ALU_SUBU 5'd2
`define ALU_SUB  5'd3
`define ALU_SLT  5'd4
`define ALU_SLTU 5'd5
`define ALU_AND  5'd6
`define ALU_OR   5'd7
`define ALU_XOR  5'd8
`define ALU_LUI  5'd9
`define ALU_SLL  5'd10
`define ALU_SRL  5'd11
`define ALU_SRA  5'd12
`define ALU_NOR  5'd13
`define ALU_MUL  5'd14
`define ALU_MULT 5'd15
`define ALU_DIV  5'd16
`define ALU_MFHI 5'd17
`define ALU_MFLO 5'd18
`define ALU_MTHI 5'd19
`define ALU_MTLO 5'd20
`define ALU_XXX  5'd31

`endif //ALUOP
