module PCAdder(
  input [31:0] A,
  input [31:0] B,
  output  [31:0] saidaAdder
);
   
    
assign  saidaAdder =(A + B);
  

endmodule
